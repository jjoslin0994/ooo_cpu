package
  

endpackage